module mesh4x4 (
    input clk,
    input reset,
    output polarity,
    input pesi_00, input [63:0] pedi_00, output peri_00, input pero_00, output [63:0] pedo_00, output peso_00,
    input pesi_01, input [63:0] pedi_01, output peri_01, input pero_01, output [63:0] pedo_01, output peso_01,
    input pesi_02, input [63:0] pedi_02, output peri_02, input pero_02, output [63:0] pedo_02, output peso_02,
    input pesi_03, input [63:0] pedi_03, output peri_03, input pero_03, output [63:0] pedo_03, output peso_03,
    input pesi_10, input [63:0] pedi_10, output peri_10, input pero_10, output [63:0] pedo_10, output peso_10,
    input pesi_11, input [63:0] pedi_11, output peri_11, input pero_11, output [63:0] pedo_11, output peso_11,
    input pesi_12, input [63:0] pedi_12, output peri_12, input pero_12, output [63:0] pedo_12, output peso_12,
    input pesi_13, input [63:0] pedi_13, output peri_13, input pero_13, output [63:0] pedo_13, output peso_13,
    input pesi_20, input [63:0] pedi_20, output peri_20, input pero_20, output [63:0] pedo_20, output peso_20,
    input pesi_21, input [63:0] pedi_21, output peri_21, input pero_21, output [63:0] pedo_21, output peso_21,
    input pesi_22, input [63:0] pedi_22, output peri_22, input pero_22, output [63:0] pedo_22, output peso_22,
    input pesi_23, input [63:0] pedi_23, output peri_23, input pero_23, output [63:0] pedo_23, output peso_23,
    input pesi_30, input [63:0] pedi_30, output peri_30, input pero_30, output [63:0] pedo_30, output peso_30,
    input pesi_31, input [63:0] pedi_31, output peri_31, input pero_31, output [63:0] pedo_31, output peso_31,
    input pesi_32, input [63:0] pedi_32, output peri_32, input pero_32, output [63:0] pedo_32, output peso_32,
    input pesi_33, input [63:0] pedi_33, output peri_33, input pero_33, output [63:0] pedo_33, output peso_33
);
    

endmodule